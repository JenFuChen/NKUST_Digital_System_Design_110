library verilog;
use verilog.vl_types.all;
entity HW3_vlg_vec_tst is
end HW3_vlg_vec_tst;
