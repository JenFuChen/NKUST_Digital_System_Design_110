library verilog;
use verilog.vl_types.all;
entity BP_tb is
end BP_tb;
