library verilog;
use verilog.vl_types.all;
entity HW3_Shoot_Darts_vlg_vec_tst is
end HW3_Shoot_Darts_vlg_vec_tst;
