library verilog;
use verilog.vl_types.all;
entity HW1_ALU_TestBench_vlg_vec_tst is
end HW1_ALU_TestBench_vlg_vec_tst;
