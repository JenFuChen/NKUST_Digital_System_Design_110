module FA(s, Carry_out, x, y, Carry_in);
input x, y, Carry_in;
output s, Carry_out;

  
endmodule

module HA(s, c, x, y);
input x, y;
output s, c;


  
endmodule

