library verilog;
use verilog.vl_types.all;
entity HW1_CSA_vlg_vec_tst is
end HW1_CSA_vlg_vec_tst;
